module mymodule

import os
import gg
import math



/**
 * Multiline comment
 * TODO   todo mark
 * FIXME  fixme mark
 *
 * "Strings" should be 'ignored' in comments
 */

// Single-line comment
// TODO FIXME
// "string" 'string'
